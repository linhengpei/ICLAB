module SMC(
    mode,
    W_0, V_GS_0, V_DS_0,
    W_1, V_GS_1, V_DS_1,
    W_2, V_GS_2, V_DS_2,
    W_3, V_GS_3, V_DS_3,
    W_4, V_GS_4, V_DS_4,
    W_5, V_GS_5, V_DS_5,   
    out_n
);
input [2:0] W_0, V_GS_0, V_DS_0;
input [2:0] W_1, V_GS_1, V_DS_1;
input [2:0] W_2, V_GS_2, V_DS_2;
input [2:0] W_3, V_GS_3, V_DS_3;
input [2:0] W_4, V_GS_4, V_DS_4;
input [2:0] W_5, V_GS_5, V_DS_5;
input [1:0] mode;

output  reg [7:0] out_n; 								
reg  [2:0]V_GS [5:0];
reg  [2:0]V_DS [5:0];
reg  [2:0]W    [5:0];

always@(*)begin  // rename
    W[0]  = W_0;
    W[1]  = W_1;
    W[2]  = W_2;
    W[3]  = W_3;
    W[4]  = W_4; 
    W[5]  = W_5;

    V_GS[0] = V_GS_0;
    V_GS[1] = V_GS_1;
    V_GS[2] = V_GS_2;
    V_GS[3] = V_GS_3;
    V_GS[4] = V_GS_4;
    V_GS[5] = V_GS_5;
    
    V_DS[0] = V_DS_0;
    V_DS[1] = V_DS_1;
    V_DS[2] = V_DS_2;
    V_DS[3] = V_DS_3;
    V_DS[4] = V_DS_4;
    V_DS[5] = V_DS_5;
end

integer i, j;
reg   Triode[5:0] ;     // Triode : 1   saturation : 0
reg  [2:0] VGS_sub1[5:0] ;     // 6 * 3 bits
reg  [3:0] VGS_sub1_2 [5:0];

always@(*)begin   // calculate  VGS_sub1  VGS_sub1_2 Triode
    for ( i = 0 ;  i <= 5 ; i = i + 1)begin 
        VGS_sub1[i] = V_GS[i] - 1;
        //VGS_sub1[i][2] = V_GS[i][2] & ( V_GS[i][1] | V_GS[i][0]);
        //VGS_sub1[i][1] = ~(V_GS[i][1] ^ V_GS[i][0]);
        //VGS_sub1[i][0] = ~V_GS[i][0];      

        VGS_sub1_2[i] = {VGS_sub1[i],1'b0};
        Triode[i] = (VGS_sub1[i] > V_DS[i]);
    end
end

reg  [2:0] Id_A [5:0];    // Id  = A * B; 
reg  [3:0] Id_B [5:0];     
reg  [2:0] Gm_A [5:0];    // Gm  = A * 2; 

always@(*)begin // calculate Id_A Id_B Gm_A
    for ( i = 0 ; i <= 5 ; i = i + 1)begin
        Id_A[i] = (Triode[i])? V_DS[i] : VGS_sub1[i] ;  
        Id_B[i] = (Triode[i])? VGS_sub1_2[i] - V_DS[i] : VGS_sub1[i] ;
        Gm_A[i] = Id_A[i]  ;
    end
end

reg  [3:0] Id_1[5:0];
reg  [3:0] Id_2[5:0];
reg  [3:0] Id_3[5:0];
reg  [7:0] Id  [5:0]; 
reg  [3:0] Gm  [5:0];
reg  [7:0] N_1 [5:0];
reg  [7:0] N_2 [5:0];
reg  [7:0] N_3 [5:0];
reg  [7:0] N   [5:0];

reg [1:0] remainder[5:0] ; 
always@(*)begin // calculate N0 ~ N5
    for (i = 0 ; i <= 5 ; i = i + 1)begin
        for (j = 0 ; j <= 3 ; j = j + 1)begin
            Id_1[i][j] = Id_A[i][0] & Id_B[i][j] ;
            Id_2[i][j] = Id_A[i][1] & Id_B[i][j] ;
            Id_3[i][j] = Id_A[i][2] & Id_B[i][j] ;
        end  
   //     Id_1[i] = (Id_A[i][0])?  Id_B[i] : 0 ;
   //     Id_2[i] = (Id_A[i][1])?  Id_B[i] : 0 ;
   //     Id_3[i] = (Id_A[i][2])?  Id_B[i] : 0 ;

       // Id[i][0] = Id_1[i][0] ;
       // Id[i][6:1] =  Id_1[i][3:1] + Id_2[i] + {Id_3[i],1'b0};
        Id[i] = Id_1[i] + {Id_2[i],1'b0} + {Id_3[i],2'b0};
        Gm[i] = {Gm_A[i],1'b0};
        N[i] = (mode[0])? Id[i] : Gm[i];
        
        // test
        /*
        case (N[i])
            1,4,7,10,13,16,19,22,25,28,31,34: remainder[i] = 1;
            2,5,8,11,14,17,20,23,26,29,32,35: remainder[i] = 2;
        endcase 

        case (N[i])
            0,1,2: N[i] = 0;
            3,4,5: N[i] = 1;
            6,7,8: N[i] = 2; 
            9,10,11: N[i] = 3; 
            12,13,14: N[i] = 4;
            15,16,17: N[i] = 5;
            18,19,20: N[i] = 6;
            21,22,23: N[i] = 7; 
            24,25,26: N[i] = 8;
            27,28,29: N[i] = 9;
            30,31,32: N[i] = 10;
            33,34,35: N[i] = 11; 
            36: N[i] = 12;
        endcase
        
        /*
        for (j = 0 ; j <= 6 ; j = j + 1)begin
            N_1[i][j] =  W[i][0] & N[i][j] ;
            N_2[i][j] =  W[i][1] & N[i][j] ;
            N_3[i][j] =  W[i][2] & N[i][j] ;
        end
        */
        N_1[i] =  (W[i][0])?   N[i] : 0 ;
        N_2[i] =  (W[i][1])?   N[i] : 0 ;
        N_3[i] =  (W[i][2])?   N[i] : 0 ;
        N[i][0] = N_1[i][0];
        N[i][7:1] = N_1[i][7:1] + N_2[i] + {N_3[i],1'b0} ;
        //N[i] = N_1[i] + {N_2[i],1'b0} + {N_3[i],2'b0} ;
        /*
        case({remainder[i],W[i]})
                5'b10010,5'b01011,5'b01100,5'b01101: N[i] = N[i] + 1; // 2 * 2 // 1 * 3 // 1 * 4
                5'b10011,5'b01110,5'b01111,5'b10100: N[i] = N[i] + 2; // 2 * 3
                5'b10101: N[i] = N[i] + 3; // 2 * 5
                5'b10110, 5'b10111: N[i] = N[i] + 4; // 2 * 6 2 * 7
        endcase
        */ 
        
        //N[i] = N[i]/3;
         
        case (N[i])
            0, 1, 2: N[i] = 0;
            3, 4, 5: N[i] = 1;
            6, 7, 8: N[i] = 2;
            9, 10, 11: N[i] = 3;
            12, 13, 14: N[i] = 4;
            15, 16, 17: N[i] = 5;
            18, 19, 20: N[i] = 6;
            21, 22, 23: N[i] = 7;
            24, 25, 26: N[i] = 8;
            27, 28, 29: N[i] = 9;
            30, 31, 32: N[i] = 10;
            33, 34, 35: N[i] = 11;
            36, 37, 38: N[i] = 12;
            39, 40, 41: N[i] = 13;
            42, 43, 44: N[i] = 14;
            45, 46, 47: N[i] = 15;
            48, 49, 50: N[i] = 16;
            51, 52, 53: N[i] = 17;
            54, 55, 56: N[i] = 18;
            57, 58, 59: N[i] = 19;
            60, 61, 62: N[i] = 20;
            63, 64, 65: N[i] = 21;
            66, 67, 68: N[i] = 22;
            69, 70, 71: N[i] = 23;
            72, 73, 74: N[i] = 24;
            75, 76, 77: N[i] = 25;
            78, 79, 80: N[i] = 26;
            81, 82, 83: N[i] = 27;
            84, 85, 86: N[i] = 28;
            87, 88, 89: N[i] = 29;
            90, 91, 92: N[i] = 30;
            93, 94, 95: N[i] = 31;
            96, 97, 98: N[i] = 32;
            99, 100, 101: N[i] = 33;
            102, 103, 104: N[i] = 34;
            105, 106, 107: N[i] = 35;
            108, 109, 110: N[i] = 36;
            111, 112, 113: N[i] = 37;
            114, 115, 116: N[i] = 38;
            117, 118, 119: N[i] = 39;
            120, 121, 122: N[i] = 40;
            123, 124, 125: N[i] = 41;
            126, 127, 128: N[i] = 42;
            129, 130, 131: N[i] = 43;
            132, 133, 134: N[i] = 44;
            135, 136, 137: N[i] = 45;
            138, 139, 140: N[i] = 46;
            141, 142, 143: N[i] = 47;
            144, 145, 146: N[i] = 48;
            147, 148, 149: N[i] = 49;
            150, 151, 152: N[i] = 50;
            153, 154, 155: N[i] = 51;
            156, 157, 158: N[i] = 52;
            159, 160, 161: N[i] = 53;
            162, 163, 164: N[i] = 54;
            165, 166, 167: N[i] = 55;
            168, 169, 170: N[i] = 56;
            171, 172, 173: N[i] = 57;
            174, 175, 176: N[i] = 58;
            177, 178, 179: N[i] = 59;
            180, 181, 182: N[i] = 60;
            183, 184, 185: N[i] = 61;
            186, 187, 188: N[i] = 62;
            189, 190, 191: N[i] = 63;
            192, 193, 194: N[i] = 64;
            195, 196, 197: N[i] = 65;
            198, 199, 200: N[i] = 66;
            201, 202, 203: N[i] = 67;
            204, 205, 206: N[i] = 68;
            207, 208, 209: N[i] = 69;
            210, 211, 212: N[i] = 70;
            213, 214, 215: N[i] = 71;
            216, 217, 218: N[i] = 72;
            219, 220, 221: N[i] = 73;
            222, 223, 224: N[i] = 74;
            225, 226, 227: N[i] = 75;
            228, 229, 230: N[i] = 76;
            231, 232, 233: N[i] = 77;
            234, 235, 236: N[i] = 78;
            237, 238, 239: N[i] = 79;
            240, 241, 242: N[i] = 80;
            243, 244, 245: N[i] = 81;
            246, 247, 248: N[i] = 82;
            249, 250, 251: N[i] = 83;
            252, 253, 254: N[i] = 84;
        endcase
            
    end
end


reg [6:0] n [5:0];
reg [6:0] temp ;
always@(*)begin // sorting N0 ~ N5 (Optimal sorting network)
    for(i = 0 ; i <= 5 ;i = i +1)
        n[i] = N[i];

    if(n[0] < n[5])begin  
        temp = n[0] ;
        n[0] = n[5] ; 
        n[5] = temp; 
    end 

    if(n[1] < n[3])begin  
        temp = n[1] ;
        n[1] = n[3] ; 
        n[3] = temp; 
    end         

    if(n[2] < n[4])begin  
        temp = n[2];  
        n[2] = n[4];
        n[4] = temp;
    end     

    if(n[1] < n[2])begin
        temp =  n[1] ;
        n[1] =  n[2] ;
        n[2] =  temp;                         
    end

    if(n[3] < n[4])begin
        temp =  n[3] ;
        n[3] =  n[4] ;
        n[4] =  temp;                         
    end

    if(n[0] < n[3])begin
        temp =  n[0] ;
        n[0] =  n[3] ;
        n[3] =  temp;                         
    end

    if(n[2] < n[5])begin  
        temp = n[2] ;
        n[2] = n[5] ; 
        n[5] = temp; 
    end         

    if(n[0] < n[1])begin
        temp =  n[0] ;
        n[0] =  n[1] ;
        n[1] =  temp;                         
    end
    
    if(n[2] < n[3])begin
        temp =  n[2] ;
        n[2] =  n[3] ;
        n[3] =  temp;                         
    end 
    
    if(n[4] < n[5])begin
        temp =  n[4] ;
        n[4] =  n[5] ;
        n[5] =  temp;                         
    end
    
    if(n[1] < n[2])begin
        temp =  n[1] ;
        n[1] =  n[2] ;
        n[2] =  temp;                         
    end

    if(n[3] < n[4])begin
        temp =  n[3] ;
        n[3] =  n[4] ;
        n[4] =  temp;                         
    end
end

reg [9:0] out_1 , out_2 , out_3 , out_4 , out_5 ;
always@(*)begin //output
    /*
    case(mode)
        2'b00:begin
                out_1 = n[3];
                out_2 = n[4];
                out_3 = n[5];
                out_n = (out_1 + out_2 +out_3);
                //out_n = (n[3] + n[4] + n[5])/3;
               end 
        2'b01:begin
                out_1 = {n[3],1'b0}  + n[3];
                out_2 = {n[4],2'b0}  ;
                out_3 = {n[5],2'b0}  + n[5];
                out_n = ((out_1 + out_2 + out_3)>>2);
                //out_n = (3 * n[3] + 4 * n[4] + 5 * n[5])/12;
               end
        2'b10:begin
                out_1 = n[0];
                out_2 = n[1];
                out_3 = n[2];
                out_n = (out_1 + out_2 +out_3);
                //out_n = (n[0] + n[1] + n[2])/3;
               end
        2'b11:begin
                out_1 = {n[0],1'b0}  + n[0];
                out_2 = {n[1],2'b0}  ;
                out_3 = {n[2],2'b0}  + n[2];
                out_n = ((out_1 + out_2 +out_3)>>2);
                //out_n = (3 * n[0] + 4 * n[1] + 5 * n[2])/12;
               end              
    endcase
    */
    out_1 = (mode[1])? n[0] : n[3] ;
    out_2 = (mode[1])? n[1] : n[4] ;
    out_3 = (mode[1])? n[2] : n[5] ;    
    out_4 = {(out_1 + out_2 + out_3),2'b0};
    
    if(mode[0])  out_5 = (out_4 + out_3 - out_1) ;  
    else         out_5 = out_4  ;
   // out_n = out_5 / 12; 
end

always@(*)begin
    out_n = 0;
    case(out_5)
        0,1,2,3,4,5,6,7,8,9,10,11  :  out_n = 0 ;
        12,13,14,15,16,17,18,19,20,21,22,23  :  out_n = 1 ;
        24,25,26,27,28,29,30,31,32,33,34,35  :  out_n = 2 ;
        36,37,38,39,40,41,42,43,44,45,46,47  :  out_n = 3 ;
        48,49,50,51,52,53,54,55,56,57,58,59  :  out_n = 4 ;
        60,61,62,63,64,65,66,67,68,69,70,71  :  out_n = 5 ;
        72,73,74,75,76,77,78,79,80,81,82,83  :  out_n = 6 ;
        84,85,86,87,88,89,90,91,92,93,94,95  :  out_n = 7 ;
        96,97,98,99,100,101,102,103,104,105,106,107  :  out_n = 8 ;
        108,109,110,111,112,113,114,115,116,117,118,119  :  out_n = 9 ;
        120,121,122,123,124,125,126,127,128,129,130,131  :  out_n = 10 ;
        132,133,134,135,136,137,138,139,140,141,142,143  :  out_n = 11 ;
        144,145,146,147,148,149,150,151,152,153,154,155  :  out_n = 12 ;
        156,157,158,159,160,161,162,163,164,165,166,167  :  out_n = 13 ;
        168,169,170,171,172,173,174,175,176,177,178,179  :  out_n = 14 ;
        180,181,182,183,184,185,186,187,188,189,190,191  :  out_n = 15 ;
        192,193,194,195,196,197,198,199,200,201,202,203  :  out_n = 16 ;
        204,205,206,207,208,209,210,211,212,213,214,215  :  out_n = 17 ;
        216,217,218,219,220,221,222,223,224,225,226,227  :  out_n = 18 ;
        228,229,230,231,232,233,234,235,236,237,238,239  :  out_n = 19 ;
        240,241,242,243,244,245,246,247,248,249,250,251  :  out_n = 20 ;
        252,253,254,255,256,257,258,259,260,261,262,263  :  out_n = 21 ;
        264,265,266,267,268,269,270,271,272,273,274,275  :  out_n = 22 ;
        276,277,278,279,280,281,282,283,284,285,286,287  :  out_n = 23 ;
        288,289,290,291,292,293,294,295,296,297,298,299  :  out_n = 24 ;
        300,301,302,303,304,305,306,307,308,309,310,311  :  out_n = 25 ;
        312,313,314,315,316,317,318,319,320,321,322,323  :  out_n = 26 ;
        324,325,326,327,328,329,330,331,332,333,334,335  :  out_n = 27 ;
        336,337,338,339,340,341,342,343,344,345,346,347  :  out_n = 28 ;
        348,349,350,351,352,353,354,355,356,357,358,359  :  out_n = 29 ;
        360,361,362,363,364,365,366,367,368,369,370,371  :  out_n = 30 ;
        372,373,374,375,376,377,378,379,380,381,382,383  :  out_n = 31 ;
        384,385,386,387,388,389,390,391,392,393,394,395  :  out_n = 32 ;
        396,397,398,399,400,401,402,403,404,405,406,407  :  out_n = 33 ;
        408,409,410,411,412,413,414,415,416,417,418,419  :  out_n = 34 ;
        420,421,422,423,424,425,426,427,428,429,430,431  :  out_n = 35 ;
        432,433,434,435,436,437,438,439,440,441,442,443  :  out_n = 36 ;
        444,445,446,447,448,449,450,451,452,453,454,455  :  out_n = 37 ;
        456,457,458,459,460,461,462,463,464,465,466,467  :  out_n = 38 ;
        468,469,470,471,472,473,474,475,476,477,478,479  :  out_n = 39 ;
        480,481,482,483,484,485,486,487,488,489,490,491  :  out_n = 40 ;
        492,493,494,495,496,497,498,499,500,501,502,503  :  out_n = 41 ;
        504,505,506,507,508,509,510,511,512,513,514,515  :  out_n = 42 ;
        516,517,518,519,520,521,522,523,524,525,526,527  :  out_n = 43 ;
        528,529,530,531,532,533,534,535,536,537,538,539  :  out_n = 44 ;
        540,541,542,543,544,545,546,547,548,549,550,551  :  out_n = 45 ;
        552,553,554,555,556,557,558,559,560,561,562,563  :  out_n = 46 ;
        564,565,566,567,568,569,570,571,572,573,574,575  :  out_n = 47 ;
        576,577,578,579,580,581,582,583,584,585,586,587  :  out_n = 48 ;
        588,589,590,591,592,593,594,595,596,597,598,599  :  out_n = 49 ;
        600,601,602,603,604,605,606,607,608,609,610,611  :  out_n = 50 ;
        612,613,614,615,616,617,618,619,620,621,622,623  :  out_n = 51 ;
        624,625,626,627,628,629,630,631,632,633,634,635  :  out_n = 52 ;
        636,637,638,639,640,641,642,643,644,645,646,647  :  out_n = 53 ;
        648,649,650,651,652,653,654,655,656,657,658,659  :  out_n = 54 ;
        660,661,662,663,664,665,666,667,668,669,670,671  :  out_n = 55 ;
        672,673,674,675,676,677,678,679,680,681,682,683  :  out_n = 56 ;
        684,685,686,687,688,689,690,691,692,693,694,695  :  out_n = 57 ;
        696,697,698,699,700,701,702,703,704,705,706,707  :  out_n = 58 ;
        708,709,710,711,712,713,714,715,716,717,718,719  :  out_n = 59 ;
        720,721,722,723,724,725,726,727,728,729,730,731  :  out_n = 60 ;
        732,733,734,735,736,737,738,739,740,741,742,743  :  out_n = 61 ;
        744,745,746,747,748,749,750,751,752,753,754,755  :  out_n = 62 ;
        756,757,758,759,760,761,762,763,764,765,766,767  :  out_n = 63 ;
        768,769,770,771,772,773,774,775,776,777,778,779  :  out_n = 64 ;
        780,781,782,783,784,785,786,787,788,789,790,791  :  out_n = 65 ;
        792,793,794,795,796,797,798,799,800,801,802,803  :  out_n = 66 ;
        804,805,806,807,808,809,810,811,812,813,814,815  :  out_n = 67 ;
        816,817,818,819,820,821,822,823,824,825,826,827  :  out_n = 68 ;
        828,829,830,831,832,833,834,835,836,837,838,839  :  out_n = 69 ;
        840,841,842,843,844,845,846,847,848,849,850,851  :  out_n = 70 ;
        852,853,854,855,856,857,858,859,860,861,862,863  :  out_n = 71 ;
        864,865,866,867,868,869,870,871,872,873,874,875  :  out_n = 72 ;
        876,877,878,879,880,881,882,883,884,885,886,887  :  out_n = 73 ;
        888,889,890,891,892,893,894,895,896,897,898,899  :  out_n = 74 ;
        900,901,902,903,904,905,906,907,908,909,910,911  :  out_n = 75 ;
        912,913,914,915,916,917,918,919,920,921,922,923  :  out_n = 76 ;
        924,925,926,927,928,929,930,931,932,933,934,935  :  out_n = 77 ;
        936,937,938,939,940,941,942,943,944,945,946,947  :  out_n = 78 ;
        948,949,950,951,952,953,954,955,956,957,958,959  :  out_n = 79 ;
        960,961,962,963,964,965,966,967,968,969,970,971  :  out_n = 80 ;
        972,973,974,975,976,977,978,979,980,981,982,983  :  out_n = 81 ;
        984,985,986,987,988,989,990,991,992,993,994,995  :  out_n = 82 ;
        996,997,998,999,1000,1001,1002,1003,1004,1005,1006,1007  :  out_n = 83 ;
        1008,1009,1010,1014,1015,1016,1017,1018,1019  :  out_n = 84 ;
        1020,1021,1022  : out_n = 85;
    endcase
end

endmodule //     37249.027464  0.01